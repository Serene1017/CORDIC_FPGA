module controller(
	);
	
endmodule
