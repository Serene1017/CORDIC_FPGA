module controller(
	output op,
	input sign,
	input comp,
	input clk
	);
	
	reg [4:0] counter;
	
	
endmodule
